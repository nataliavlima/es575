library verilog;
use verilog.vl_types.all;
entity Exp2b_vlg_sample_tst is
    port(
        v0              : in     vl_logic;
        v1              : in     vl_logic;
        v2              : in     vl_logic;
        v3              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Exp2b_vlg_sample_tst;
