library verilog;
use verilog.vl_types.all;
entity Exp2b_vlg_vec_tst is
end Exp2b_vlg_vec_tst;
